`timescale 1ns/1ps

module top (
    // 16MHz clock
    input CLK,

    // USB pull-up resistor
    output USBPU,

    // GPIO Inputs.
    input PIN_1,
    input PIN_2,
    input PIN_3,
    input PIN_4,
    input PIN_5,
    input PIN_6,
    input PIN_7,
    input PIN_8,
    input PIN_9,
    input PIN_10,
    input PIN_11,
    input PIN_12,
    input PIN_13,
    input PIN_14,
    input PIN_15,

    input PIN_16,

    // GPIO Outputs.
    inout PIN_17,
    inout PIN_18,
    inout PIN_19,
    inout PIN_20,
    inout PIN_21,
    inout PIN_22,
    inout PIN_23,
    inout PIN_24
);

    // drive USB pull-up resistor to '0' to disable USB
    assign USBPU = 0;

    // External flag to turn output on.  Usually a chip enable signal.
    wire output_on;
    assign output_on = PIN_16;

    // Address inputs.
    wire a0;
    wire a1;
    wire a2;
    wire a3;
    wire a4;
    wire a5;
    wire a6;
    wire a7;
    wire a8;
    wire a9;
    wire a10;
    wire a11;
    wire a12;
    wire a13;
    wire a14;

    assign a0 = PIN_1;
    assign a1 = PIN_2;
    assign a2 = PIN_3;
    assign a3 = PIN_4;
    assign a4 = PIN_5;
    assign a5 = PIN_6;
    assign a6 = PIN_7;
    assign a7 = PIN_8;
    assign a8 = PIN_9;
    assign a9 = PIN_10;
    assign a10 = PIN_11;
    assign a11 = PIN_12;
    assign a12 = PIN_13;
    assign a13 = PIN_14;
    assign a14 = PIN_15;

    wire [10:0] rom_address;
    assign rom_address = {1'b0, 1'b0, a8, a7, a6, a5, a4, a3, a2, a1, a0};
    wire [5:0] rom_select;
    assign rom_select = {a14, a13, a12, a11, a10, a9};

    // Data output.
    reg data0;
    reg data1;
    reg data2;
    reg data3;
    reg data4;
    reg data5;
    reg data6;
    reg data7;

    // Allow for high impedance mode in data lines.
    wire data0tri;
    assign data0tri = (!output_on) ? data0 : 1'bZ;
    wire data1tri;
    assign data1tri = (!output_on) ? data1 : 1'bZ;
    wire data2tri;
    assign data2tri = (!output_on) ? data2 : 1'bZ;
    wire data3tri;
    assign data3tri = (!output_on) ? data3 : 1'bZ;
    wire data4tri;
    assign data4tri = (!output_on) ? data4 : 1'bZ;
    wire data5tri;
    assign data5tri = (!output_on) ? data5 : 1'bZ;
    wire data6tri;
    assign data6tri = (!output_on) ? data6 : 1'bZ;
    wire data7tri;
    assign data7tri = (!output_on) ? data7 : 1'bZ;

    assign PIN_17 = data0tri;
    assign PIN_18 = data1tri;
    assign PIN_19 = data2tri;
    assign PIN_20 = data3tri;
    assign PIN_21 = data4tri;
    assign PIN_22 = data5tri;
    assign PIN_23 = data6tri;
    assign PIN_24 = data7tri;

    wire [15:0] memory_data_out_0;
    wire [15:0] memory_data_out_1;
    wire [15:0] memory_data_out_2;
    wire [15:0] memory_data_out_3;
    wire [15:0] memory_data_out_4;
    wire [15:0] memory_data_out_5;
    wire [15:0] memory_data_out_6;
    wire [15:0] memory_data_out_7;
    wire [15:0] memory_data_out_8;
    wire [15:0] memory_data_out_9;
    wire [15:0] memory_data_out_10;
    wire [15:0] memory_data_out_11;
    wire [15:0] memory_data_out_12;
    wire [15:0] memory_data_out_13;
    wire [15:0] memory_data_out_14;
    wire [15:0] memory_data_out_15;
    wire [15:0] memory_data_out_16;
    wire [15:0] memory_data_out_17;
    wire [15:0] memory_data_out_18;
    wire [15:0] memory_data_out_19;
    wire [15:0] memory_data_out_20;
    wire [15:0] memory_data_out_21;
    wire [15:0] memory_data_out_22;
    wire [15:0] memory_data_out_23;

    initial begin
    end

    always @(posedge clk_40mhz) begin
      if (rom_select == 0) begin
            data7 <= memory_data_out_0[14];
            data6 <= memory_data_out_0[12];
            data5 <= memory_data_out_0[10];
            data4 <= memory_data_out_0[8];
            data3 <= memory_data_out_0[6];
            data2 <= memory_data_out_0[4];
            data1 <= memory_data_out_0[2];
            data0 <= memory_data_out_0[0];
      end else if (rom_select == 1) begin
            data7 <= memory_data_out_1[14];
            data6 <= memory_data_out_1[12];
            data5 <= memory_data_out_1[10];
            data4 <= memory_data_out_1[8];
            data3 <= memory_data_out_1[6];
            data2 <= memory_data_out_1[4];
            data1 <= memory_data_out_1[2];
            data0 <= memory_data_out_1[0];
      end else if (rom_select == 2) begin
            data7 <= memory_data_out_2[14];
            data6 <= memory_data_out_2[12];
            data5 <= memory_data_out_2[10];
            data4 <= memory_data_out_2[8];
            data3 <= memory_data_out_2[6];
            data2 <= memory_data_out_2[4];
            data1 <= memory_data_out_2[2];
            data0 <= memory_data_out_2[0];
      end else if (rom_select == 3) begin
            data7 <= memory_data_out_3[14];
            data6 <= memory_data_out_3[12];
            data5 <= memory_data_out_3[10];
            data4 <= memory_data_out_3[8];
            data3 <= memory_data_out_3[6];
            data2 <= memory_data_out_3[4];
            data1 <= memory_data_out_3[2];
            data0 <= memory_data_out_3[0];
      end else if (rom_select == 4) begin
            data7 <= memory_data_out_4[14];
            data6 <= memory_data_out_4[12];
            data5 <= memory_data_out_4[10];
            data4 <= memory_data_out_4[8];
            data3 <= memory_data_out_4[6];
            data2 <= memory_data_out_4[4];
            data1 <= memory_data_out_4[2];
            data0 <= memory_data_out_4[0];
      end else if (rom_select == 5) begin
            data7 <= memory_data_out_5[14];
            data6 <= memory_data_out_5[12];
            data5 <= memory_data_out_5[10];
            data4 <= memory_data_out_5[8];
            data3 <= memory_data_out_5[6];
            data2 <= memory_data_out_5[4];
            data1 <= memory_data_out_5[2];
            data0 <= memory_data_out_5[0];
      end else if (rom_select == 6) begin
            data7 <= memory_data_out_6[14];
            data6 <= memory_data_out_6[12];
            data5 <= memory_data_out_6[10];
            data4 <= memory_data_out_6[8];
            data3 <= memory_data_out_6[6];
            data2 <= memory_data_out_6[4];
            data1 <= memory_data_out_6[2];
            data0 <= memory_data_out_6[0];
      end else if (rom_select == 7) begin
            data7 <= memory_data_out_7[14];
            data6 <= memory_data_out_7[12];
            data5 <= memory_data_out_7[10];
            data4 <= memory_data_out_7[8];
            data3 <= memory_data_out_7[6];
            data2 <= memory_data_out_7[4];
            data1 <= memory_data_out_7[2];
            data0 <= memory_data_out_7[0];
      end else if (rom_select == 8) begin
            data7 <= memory_data_out_8[14];
            data6 <= memory_data_out_8[12];
            data5 <= memory_data_out_8[10];
            data4 <= memory_data_out_8[8];
            data3 <= memory_data_out_8[6];
            data2 <= memory_data_out_8[4];
            data1 <= memory_data_out_8[2];
            data0 <= memory_data_out_8[0];
      end else if (rom_select == 9) begin
            data7 <= memory_data_out_9[14];
            data6 <= memory_data_out_9[12];
            data5 <= memory_data_out_9[10];
            data4 <= memory_data_out_9[8];
            data3 <= memory_data_out_9[6];
            data2 <= memory_data_out_9[4];
            data1 <= memory_data_out_9[2];
            data0 <= memory_data_out_9[0];
      end else if (rom_select == 10) begin
            data7 <= memory_data_out_10[14];
            data6 <= memory_data_out_10[12];
            data5 <= memory_data_out_10[10];
            data4 <= memory_data_out_10[8];
            data3 <= memory_data_out_10[6];
            data2 <= memory_data_out_10[4];
            data1 <= memory_data_out_10[2];
            data0 <= memory_data_out_10[0];
      end else if (rom_select == 11) begin
            data7 <= memory_data_out_11[14];
            data6 <= memory_data_out_11[12];
            data5 <= memory_data_out_11[10];
            data4 <= memory_data_out_11[8];
            data3 <= memory_data_out_11[6];
            data2 <= memory_data_out_11[4];
            data1 <= memory_data_out_11[2];
            data0 <= memory_data_out_11[0];
      end else if (rom_select == 12) begin
            data7 <= memory_data_out_12[14];
            data6 <= memory_data_out_12[12];
            data5 <= memory_data_out_12[10];
            data4 <= memory_data_out_12[8];
            data3 <= memory_data_out_12[6];
            data2 <= memory_data_out_12[4];
            data1 <= memory_data_out_12[2];
            data0 <= memory_data_out_12[0];
      end else if (rom_select == 13) begin
            data7 <= memory_data_out_13[14];
            data6 <= memory_data_out_13[12];
            data5 <= memory_data_out_13[10];
            data4 <= memory_data_out_13[8];
            data3 <= memory_data_out_13[6];
            data2 <= memory_data_out_13[4];
            data1 <= memory_data_out_13[2];
            data0 <= memory_data_out_13[0];
      end else if (rom_select == 14) begin
            data7 <= memory_data_out_14[14];
            data6 <= memory_data_out_14[12];
            data5 <= memory_data_out_14[10];
            data4 <= memory_data_out_14[8];
            data3 <= memory_data_out_14[6];
            data2 <= memory_data_out_14[4];
            data1 <= memory_data_out_14[2];
            data0 <= memory_data_out_14[0];
      end else if (rom_select == 15) begin
            data7 <= memory_data_out_15[14];
            data6 <= memory_data_out_15[12];
            data5 <= memory_data_out_15[10];
            data4 <= memory_data_out_15[8];
            data3 <= memory_data_out_15[6];
            data2 <= memory_data_out_15[4];
            data1 <= memory_data_out_15[2];
            data0 <= memory_data_out_15[0];
      end else if (rom_select == 16) begin
            data7 <= memory_data_out_16[14];
            data6 <= memory_data_out_16[12];
            data5 <= memory_data_out_16[10];
            data4 <= memory_data_out_16[8];
            data3 <= memory_data_out_16[6];
            data2 <= memory_data_out_16[4];
            data1 <= memory_data_out_16[2];
            data0 <= memory_data_out_16[0];
      end else if (rom_select == 17) begin
            data7 <= memory_data_out_17[14];
            data6 <= memory_data_out_17[12];
            data5 <= memory_data_out_17[10];
            data4 <= memory_data_out_17[8];
            data3 <= memory_data_out_17[6];
            data2 <= memory_data_out_17[4];
            data1 <= memory_data_out_17[2];
            data0 <= memory_data_out_17[0];
      end else if (rom_select == 18) begin
            data7 <= memory_data_out_18[14];
            data6 <= memory_data_out_18[12];
            data5 <= memory_data_out_18[10];
            data4 <= memory_data_out_18[8];
            data3 <= memory_data_out_18[6];
            data2 <= memory_data_out_18[4];
            data1 <= memory_data_out_18[2];
            data0 <= memory_data_out_18[0];
      end else if (rom_select == 19) begin
            data7 <= memory_data_out_19[14];
            data6 <= memory_data_out_19[12];
            data5 <= memory_data_out_19[10];
            data4 <= memory_data_out_19[8];
            data3 <= memory_data_out_19[6];
            data2 <= memory_data_out_19[4];
            data1 <= memory_data_out_19[2];
            data0 <= memory_data_out_19[0];
      end else if (rom_select == 20) begin
            data7 <= memory_data_out_20[14];
            data6 <= memory_data_out_20[12];
            data5 <= memory_data_out_20[10];
            data4 <= memory_data_out_20[8];
            data3 <= memory_data_out_20[6];
            data2 <= memory_data_out_20[4];
            data1 <= memory_data_out_20[2];
            data0 <= memory_data_out_20[0];
      end else if (rom_select == 21) begin
            data7 <= memory_data_out_21[14];
            data6 <= memory_data_out_21[12];
            data5 <= memory_data_out_21[10];
            data4 <= memory_data_out_21[8];
            data3 <= memory_data_out_21[6];
            data2 <= memory_data_out_21[4];
            data1 <= memory_data_out_21[2];
            data0 <= memory_data_out_21[0];
      end else if (rom_select == 22) begin
            data7 <= memory_data_out_22[14];
            data6 <= memory_data_out_22[12];
            data5 <= memory_data_out_22[10];
            data4 <= memory_data_out_22[8];
            data3 <= memory_data_out_22[6];
            data2 <= memory_data_out_22[4];
            data1 <= memory_data_out_22[2];
            data0 <= memory_data_out_22[0];
      end else if (rom_select == 23) begin
            data7 <= memory_data_out_23[14];
            data6 <= memory_data_out_23[12];
            data5 <= memory_data_out_23[10];
            data4 <= memory_data_out_23[8];
            data3 <= memory_data_out_23[6];
            data2 <= memory_data_out_23[4];
            data1 <= memory_data_out_23[2];
            data0 <= memory_data_out_23[0];
      end else if (rom_select == 63) begin
        // 6502 reset and interrupt vectors.
        if (rom_address == 506) begin // Low byte NMI interrupt.
          data7 <= 0;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end else if (rom_address == 507) begin // High byte NMI interrupt.
          data7 <= 0;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end else if (rom_address == 508) begin // Low byte reset vector.
          data7 <= 0;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end else if (rom_address == 509) begin // High byte reset vector.
          data7 <= 1;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end else if (rom_address == 510) begin // Low byte interrupt.
          data7 <= 0;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end else if (rom_address == 511) begin // High byte interrupt.
          data7 <= 0;
          data6 <= 0;
          data5 <= 0;
          data4 <= 0;
          data3 <= 0;
          data2 <= 0;
          data1 <= 0;
          data0 <= 0;
        end
      end
    end

    // Create a 40MHz clock.
    wire clk_40mhz;
    SB_PLL40_CORE #(
      .DIVR(0),
      .DIVF(39),
      .DIVQ(4),
      .FILTER_RANGE(3'b001),
      .FEEDBACK_PATH("SIMPLE"),
      .DELAY_ADJUSTMENT_MODE_FEEDBACK("FIXED"),
      .FDA_FEEDBACK(4'b0000),
      .DELAY_ADJUSTMENT_MODE_RELATIVE("FIXED"),
      .FDA_RELATIVE(4'b0000),
      .SHIFTREG_DIV_MODE(2'b00),
      .PLLOUT_SELECT("GENCLK"),
      .ENABLE_ICEGATE(1'b0)
    ) pll (
      .REFERENCECLK(CLK),
      .PLLOUTCORE(clk_40mhz),
      .RESETB(1'b1),
      .BYPASS(1'b0)
    );

    ////
    // Insert BRAM definitions after this point.
    ////

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0011111111111111010101010000010111000000111100110111111111111111110011001100001100111111111111111111111100000110110000001111001101010101011101011100110001100011001111111111111111111111010101001100000011110011000101010111011111001100011000110001010101100010),
      .INIT_1(256'b0110110001000001001111111111111111111100010101101100000011110011101111111111111111001100110000110011110101010101011111111010101111101000010100111000000010100010010001000100000110011101110101110111110100000000010000101101000100101000000000000110110011000001),
      .INIT_2(256'b1100010001001001011010100010010101100100111000010010011000000010010000000100000011010111101001110000010000101000100111010111011101010100100000011110001001010001000000000000001011100100110000110001010101110101110111000010110101000000011100111101110101110111),
      .INIT_3(256'b0101010110000001111000100101000100000000000110101110010010010011100101010101110101111111001000000110000011110001001000100001100101000100000100011000001010110011010000000011100110001000001000110100010011000001101000100001000001000000000110011010000010000011),
      .INIT_4(256'b0101010100000000110101111111011101010000011010011100100100100111000000001100000011100111010100010100000001100100111001011001011110010000010110000110101000100000001100001110010000100110000010100000000000000000110001101010011000010001011010001001110101110111),
      .INIT_5(256'b1000000000011000011110110010000000100000111100010111001001100011010000000001010011000110101100100000010000101000100111000010001001000000100000001011001001000100000100000111001011110100110000101100000000001000001111100011000000100100101000000010001000110101),
      .INIT_6(256'b0000000010010000111100100001010000010101011111111010000010000010110000000101100100101110001000000110010011100001001001110011100101010001000000001000001011100010010100000110100110011000011000100100000010000001101000110000000000010000011110001011000011000010),
      .INIT_7(256'b0000000000010000110000101011001100000101001010001100110001100011000000001100000111110111000000000000000010000001111100001100001110000000000110010110111000110001001000011010000101110011001010100000000000000000110100101110001100000000001110001100110000110011),
      .INIT_8(256'b1101010100001000011010100111000100100000101100010110011010010011000101010101010110000010101000100100000001111001100011000010001001000100110000011010001000010000010101001001011011100000100000101100000000011101001110100111000000100000101100010111001010010100),
      .INIT_9(256'b0000000011000101111100100100000101000000100010111010000110000010100100000101100000111111011101010010000010100000011000101101100100010101010101011100011011100011000101010111110111011101001000110100000011010001101000100001000001000100100110011011010111010111),
      .INIT_A(256'b0100000100000001110100101110001100010100001011001101110100100010010000001000000011110010010000010001010010110100111101011000001010000001000010010111101001100001001101001110010001110111100010100000000001010100110100101110001100010100011111001100100100100010),
      .INIT_B(256'b1000010000001000011011100110000100100100111100010111001110100010000000000101000111010010111000110001000100111100110111010010001001010101110101011111001001000001000100011110011011110101100000101100000100001101011110100110000100110001111101000111011110100000),
      .INIT_C(256'b0000010010000000101000100100010001010001101010101010000111010011110100000100100100101010001100010110010010110001001000101011100101010100000101001000001010110010010000000011100110001000001000110100010011000001101101110101010100000000101010001110000011010011),
      .INIT_D(256'b0000000000010000110001101011001100010101011111011101110100100010010000001101000110100010000100010100011000010001101000001001001111000000000110010010101101110000011001001110000101100010101110100100000001010000100001101010001001000000001011001001110100110011),
      .INIT_E(256'b1000000000011100011010100011000100110101111101010010100000000010010000000101000111000010101000110000000100101000100110000111001000010101110101011010001000000000010000100101001110110101110101111100010001001001001111110111010101110101101000010110100001010001),
      .INIT_F(256'b0101010010010100101000100001000001000010000110111010000010000011110001000100100100101010001101000111000110100000001010000001100001010000000100011000011110100011010001000110100110001000001100100101010010010100111000100000000100000110000010001010010010000010)
    ) ram0 (
      .RDATA(memory_data_out_0),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1000100000001000111010110111101110100010000101001110010010011001001000101110100001010001000000001000001110110010011100101110101101000000000001001001111110110010000110100101000010011100000011011010101000101010111000110101000110100000100111000110011010110011),
      .INIT_1(256'b1100001010100110001111010001001000010000010100001001111010110011000010100000000011001001010110011010101000111110111001100001000110100000110010000111001110101010000000010001000111010010111000110110100000000100000101010001000010011010111100100001111000010000),
      .INIT_2(256'b1010101001101010111100110000000010100001100111010111100001000011010000000000010010010111101100100011100001011000000101000001010010001010101000100100101101010001100010000001110011101110001110111010001001000000111100011000100000101001000101000101000001000001),
      .INIT_3(256'b0010100000100000010000010101000110001010101101100100111000010001100010000100100011111011001010101010001101000000111100001100100101101000000011000001010100010000100100101111001000111100000111110000000000000000110010111111001100001010000101001100110000011001),
      .INIT_4(256'b1110001000000100101101011001100000111000011100000001010001000001100000101010001001101001011100110000000000010100110011101011001100001010010000001101100100001000101010110110101111110010010000011110000010001100001111010001101000010000010100001001011011100010),
      .INIT_5(256'b0000000001000000110110111010001000001011010001011101100001001001111010100010111010110111000100001011000011011000001111000110011000000000000000001100001111110011001010000011110001000100000100011000101011100010010110110000000010001001010011001111101001101011),
      .INIT_6(256'b1010000010001000011010010111101100000000000101001100011010110011001010001100000001010001000000001000101111110010010110100100000111001000000011001011111100111010101100100101000010110100110011010010100000101000010000010101000110000010101101100110110000111011),
      .INIT_7(256'b1101111110110111010110110000000011011000010011001011101100101011101000100000000011100001110110010011100110000100000000000000000011000111111100110010110110000010010001000000010010011110101000100100101000000100100111010001100010111010011110101011011001010000),
      .INIT_8(256'b0011100110011000000000000000000011000111111100110010110110001010010001000000010011011111101101110101101100000000110110000100110010111011001011101010001000000000111000011101100100111001100001110000000000000000110001111111001100101101100010000100010000000100),
      .INIT_9(256'b0101100100000000110110001100011010111011001110101010001000000000111000011101100100111001100110110000000000000000110001111111001100101101101000000100010000000100110111111011011101011011000000001101100001001100101110110010111110100010000000001110000111011001),
      .INIT_A(256'b0010001000000010010001010101000110000111101000100100111000000100110111010001110101011001000000001101100011000110001110010001000110101010100010001110001101010001101100011001110000101000101000000100010101010001100001111010001001001110000001001101110100011101),
      .INIT_B(256'b0111001001001110000100010001010110000010101000100100101101010001100110010100100010101010100010001110011101010001101001011000100001100110000011000101010100010101110100111010001001011010010001001001100100011100101010101000100011100011010100011011000110011101),
      .INIT_C(256'b0110011101110011000001010000000011000110101001100101111100010101110110010000100011111010110011001011001101000000101000001000100001100011011100010001000101000001100000101010001001001111010100011000110100001000111011101000110011110111000101011111000110001000),
      .INIT_D(256'b0011001101101110000000000000000011000011111100110001101101000101100010000000100011101111110110011010011100000000111001001000110001110111001111010101000100000000110100101110011000011011010000011000100000001000111010111101100110110011010001001010000010001000),
      .INIT_E(256'b0010011110000010010001000000010011010111101101110101101100000000110110000100110010111011110011011010001000000000111000011101100100110011110100000000000000000000110001111111001100001111000000001100110000001100111111111001110111110011000000001111000011001100),
      .INIT_F(256'b0010001010001010010000010101000110010011111101100000101000000000110011010101100110101111100010001110011000000100111101011001110101110011100010000101000001000100100100111111001000001010000000001100100101011001101110111101100110100010000000001110010111011001)
    ) ram1 (
      .RDATA(memory_data_out_1),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1011001101010001101000001000100001101011111110110000010100000000110001001010011001110111011011100101000100000000110110101110011000111011111110101010101000000010110000011111100100001111000000001100110000001100011111111110111011111011000000001101000011100110),
      .INIT_1(256'b0001000101010101100000001010001001100011110100010000010100000000110011101010011001111111111011101111101100000010110100001110110000011011010101001000100000001000011010111111101110101111000000001100010010100110010101011100010011011001100000101111101001100100),
      .INIT_2(256'b0001010000000001100010101010001001101011111110111010111100000010110001001010110001011111010001001101100100001000011110101110111010111110000000001000000010100010010000011101001110001101100000101110111000100100111101110100010011110001100010000111101011101110),
      .INIT_3(256'b1011111000000111100000001010100001001011010100011000110100001000011011101010111011111111010001001101000110100010010100001100110010011100100001101010101000100000111000110101000110100101100010000110111010101110010101010100010011010001101000100111001011000110),
      .INIT_4(256'b1001110000011001001010101010101011101011010100011000010110100010010001001000111011011101110001101111101100100000111100100100010010110100100110000010101010101010010000010101000110000101101000100110011010001100010101010100010011011011101000100111101011101110),
      .INIT_5(256'b1001010010110111000000001010000011001001110100111010111100100000111001100000010011110101110011000111101110101010010100000100010010010100101101100010001010001010010000010101000110001111101000100110111010101110111111110100011011010001101010000101101001000100),
      .INIT_6(256'b1011111001100001101000100000000011100001110110010010111110101010010001000000010011010101111001100111001110100000010100000100010010011110111000100010101010101010111010110101001110000101101010000100111000000100110111010100110001111011101010101111101001000100),
      .INIT_7(256'b0011111011101111000000000000000011000001111100110010011110100010010001000000010011011111111001100111101110101010111110100100011010010100111011000000101000000000110010010101100100101111101010101110111000000100110101011110011001010001101000101101100011000110),
      .INIT_8(256'b0111011110101000010000000101000110001010101000110110111011101011101111100000001011010101111011000101101100000000110110000100110000111110111110101010101000000000110000011111001100000101101010001100110010000110111111110110010011110011000000001111000011001100),
      .INIT_9(256'b0110111011101011111111110001001011010001101010000101101001000100100111010101110100101010101010101110101001010001100100011010001100000000101010101100110111010011101111110111010111110111000000011110000011011100001011111010101001000100000001001001010111110111),
      .INIT_A(256'b0101101001000100100111010101110100101010101010101110101001010001100100011010011000000010000000001100110111010011101111110111010111110111000000011110000011011100001011111010101001000100000001001001010111110111011101111010101001000000010100011000101010100110),
      .INIT_B(256'b1110101001010001100100011010011100000010000000101100110111010011101111110111010111110111000000011110000011011100001011111010101001000100000001001001010111110111011111010000000001000000010100011000101010100111011011101110101111111111000100101101000110101000),
      .INIT_C(256'b1100110111010011101111110111010111110111000000011110000011011100001011111010101001000100000001001001010111110111011111010000001001000000010100011000101010110010011011101110101111111111000100101101000110101000010110100100010010011101010111010010101010101010),
      .INIT_D(256'b1110000011011100001011111010101001000100000001001001010111110111011111010000100001000000010100011000101010110011011011101110101111111111000100101101000110101000010110100100010010011101010111010010101010101010111010100101000110010001101100100000001000001000),
      .INIT_E(256'b1001010111110111011111010000101001000000010100011000101010110110011011101110101111111111000100101101000110101000010110100100010010011101010111010010101010101010111010100101000110010001101100110000001000001010110011011101001110111111011101011111011100000001),
      .INIT_F(256'b1000101010110111011011101110101111111111000100101101000110101000010110100100010010011101010111010010101010101010111010100101000110010001101101100000001000100000110011011101001110111111011101011111011100000001111000001101110000101111101010100100010000000100)
    ) ram2 (
      .RDATA(memory_data_out_2),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0100001001010100100011011000001001101100000001000001010101011101110111011000001001101000010100010010100110010001111011101100101111111111000100001101000100101010110100001110110000011101010101011010001010001000110010001101100100011100000100001010100010000010),
      .INIT_1(256'b0001010101011101110101010010001001000000010110010010000110010110010001000100100111011101001100101101000100101010010110100110111000110101111101010000000000001000110000000111001100010100000110010000000000100010010001011101000110011101110101110101110110100001),
      .INIT_2(256'b0000000100011101110011000110001111010101001110100101101100101010011100001110010010010101110101010000000000101010010010000101000100010100000111101000100000100010110001010111101100011111011111110111010110100001110000001101011000000101100010000100110000000100),
      .INIT_3(256'b1111101100000000111110100100010010110101110101111000000010000000110000100101100100011100000101010010100000000000010001010101000110011101110101111101010110000011010000001101110000001101000000000100010000001100100101010111011101010101001000000110000011010011),
      .INIT_4(256'b1010000010000010111010101101000100010110010000001010000010001000010001011101100110111111010101011101010100101011011000101101110010100111101000100100010000001110100111010101110111110101101000001110101001010001000000110110000011100100110000110101110100010010),
      .INIT_5(256'b0010100010001000010011010101000100111111111101010101011100001001011000001101110000101111101010000110110000000100100101010111111101110111101010001100101011110011001010010100000111000100010000010101010110010010010100010000100001011010010001000001111111111111),
      .INIT_6(256'b1111010110000011110000001101010010000111000010000100110000000100100101010111111101011111001010100110000011110001000000011110110011100110010000010101011100011000111100011000001011010000110001001001011101011101000010000000000001000000111110110001010001000001),
      .INIT_7(256'b1100110010000110100111111101010111110111000000000100001001010011101000011100011101000100011010111111111100010000010100110010000011110000110001100001010111111101101010100000000001100010110100111011010011000110000000100000100011101111010100010001011101011101),
      .INIT_8(256'b0100000001011001100010010111001011000100011010110101111100111010011100011010000001010000010011001001010101110111000000000000100001001000011100111011110011101111100010001000001001001101111100011011111101111111110111011000001101101000010101000000011100001010),
      .INIT_9(256'b1101011100011000010110010000000001010000011011101001110101011101001010000000000001000000010100111001010011010010000000000000100011001101011100111001010111010111010101011000100101001000010101000000010100001000110001000010011000010101010101110111010110000010),
      .INIT_A(256'b0101011100000000111000001001110101000100001101011010111000000000110000000110101011001011100011001010011010100010010101011110110111011001000010000110100000010101010000100101010010001100100000101110101011001000111101110000010110100100100010001001010010000000),
      .INIT_B(256'b0010101000101110010001100011000100100010110100110000001100001000001101111101010011010000010010111000000100101011101001011000001000111110111000010101000001000001100010010011001111011101100010000001010111001000110100001100100101101100010001001111111111000000),
      .INIT_C(256'b0101010110101000100000010010101001000000111010011000000000101110010011001011100111000000001111100101000110011011000100000101000011101110111011101011111111111101101011001110100111001000110011001010101011011001111111110000000010101000000001001110100001000011),
      .INIT_D(256'b0100101001111111110100000110101101001010011010111000010100101010010011110111101110000000011111110111110110100000100000000110101001001010110010011000000000101110110001101011000111000100011011100100001010001000100000000110101101000010010001101000000000111010),
      .INIT_E(256'b1110110001001100110001011110011011110101101010100100100011000011001011111010101011101101010110011100100010110111000000000010011110011000010110001100010011000100010100000010011111010101100000000000000101110111100001000110101101001101011111011101010100101010),
      .INIT_F(256'b0000010101000000100010001001001011000101100000001011110101000101010110000100000110101010011010001110001100000000101101001000100101010000110000111110101001000100001010101111101111111101000000000000100010110000010000100100000110001000100001100110111010111011)
    ) ram3 (
      .RDATA(memory_data_out_3),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0001110101010101110101001000000001000100011110110000100000000101111010001011001110011001110001101111100111100110101000100000000011001000100110011111010110010010110001001100000110010110000010000100100001000000111111100010000010100110000000001011111010001000),
      .INIT_1(256'b0100011001000001100111011101011101111100000001001100000011010001000001010010101000001000010000010001010101111111010111001000011001000100010110011001110101110111111111100010000011100010010100011010111010001000101000001100001111010100110101011000011001001001),
      .INIT_2(256'b0011110101010101010111000000000001001000110100110111101011111111101011000100000110011101111101111111111010001010111001100101000100101010111010101110110000000100000010001010000011101110100000101111111101010001011110111010101010101101010001000000100110100000),
      .INIT_3(256'b1100010011111011001010000100010101000101100000101000000000100000100101000011110011000000110000011000000111011100000001000000000010010101111101011101010000001100110000000101001111010100010111111000010001100011100101010111111111010100100001100100010001010001),
      .INIT_4(256'b1100100001010011000011100000100000101010011010110011110101010111011111100000101001101110110110010100000001000000000100010000010100010000010100000001111101010111011111100000001001000000010100011111100101010101000001000100000110011101010101010101010000001010),
      .INIT_5(256'b1101110000001010010011100111001100101010010011010111101100100000001010000010100100101110011010010100100101000000010101000000010011011001000010000101101001001110010010100110000100101001011101100010110000100000011110101100000000111101010111110101010000001000),
      .INIT_6(256'b0101010000000000010010101101000101011011011111110010111001100011001111011101110101111100101000100100010001010001010000000100000000010101000000010001101001111000001111111101011101111100001010100110100011010001001011000000100000101000111010010001010101010101),
      .INIT_7(256'b0000000101010100000011001010001001111111010001000001111111001110001111011111010101011100101011100100100011111001010100000101010100000100010000010001111111010111010111100000010001101100111110110110100011000011001010011101111000001100101000000001010101010101),
      .INIT_8(256'b0000010000000000010101010101010001100110111000010100000001000000011101101010001000010000111100100101010101000001010101010000000000000001000000000000010001000001000111111111011101110110100010100100010001010001000111010010101001010001000000000100000001000001),
      .INIT_9(256'b0101010000000100010001000101000100000000010000000100111000101110000010100010000001001100101010100000101000000011010000000001000100000000000000000100000010010001000000000000000001000100010000010001000101000100010100010100010001000000010000000000000000010101),
      .INIT_A(256'b0001010101010101110101001010001001001110110100110101110111001001010110011010001000011111010111110101110010001010100001001101101000000001000000000100011011001011000111111101010101011110001011000100101001110011010110100101110100001100111010010001111101010101),
      .INIT_B(256'b1111000110101010011110101110110001010000110000101010000000100001101000010010100010100000100000001011010010011100000000000000000111110000111000011110000001001001101000010101011010100100000010101111010100100110111100010010101010100100100000100000010001000001),
      .INIT_C(256'b1111110100000010001000000000000100100110011010110010000000000011001100100001101101110111110011000001010101000100010000010100000000000000000000010101110000010110001000100000011001010101000000001110100001000001000000010101010010001100000000000101010100001111),
      .INIT_D(256'b1011110000001010000010000010001001100110000110010110001001100000011101000010100000100110001010000100110101000000010101010000000010101000000010000100110000011011010011010011010101110101001000100110000001100001001000111101010000100100000010100100010101011000),
      .INIT_E(256'b0100000001010001000010011000100000001000011010010111001001110111001001001100100100110101111101110101010000000100010001000101000100010101010101010111011010101000011000101101001101110100011111110010010011000001001101010101110101110100101010000100010001010001),
      .INIT_F(256'b0101000001000001011000101110101001100011000001000000111010001000011000001110000000001010101111110000111010101000010101010101010101000100010000010000100010000100010010001001001100100000101011100110010011000011001101001000101000011111111101010101010000000100)
    ) ram4 (
      .RDATA(memory_data_out_4),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1000100010100010000010001000100010010101011100101000000010001000100111110111001110001000111100111000000010101000101000000010001000001000000000000000100000101010100001000110011110110101011011111000000000100010000011000000111010001000001000100000100000101000),
      .INIT_1(256'b1000101010101000100000000010100000000000000000001100100100011101111000010001000010000100011101110100101100000001100010001000001010100000000000101000000001100010100000000000000010001000100000100000100010001010100000000010001010000000100010001000101000101000),
      .INIT_2(256'b0011100001110010110100000101101111000001110010110000110001100100001001001111000111000001100011110000111001000101010110000100010110000000101000100000101101101111010010010100000011100011100101001100001110011001111000011000110010110101010111011100000100101000),
      .INIT_3(256'b0010001100000100100110101111001001100000100000001001010010011000001100100101001011001010101000101001100111001001000100001101100001000000111001001101011101000101000100001101000011100000110001100110111110011111100110100101000001001010000000001011000010000110),
      .INIT_4(256'b1100011100100011001111001000000011110000000001101100001100000011010100000000010111001010001101100010000010010001111000010000001011011010000001111100100010011100101001000000001000101000001000100010000000000000000000011100010100100000110000001100000010001001),
      .INIT_5(256'b1100000011011000100011110110011111101000111100100001111110000001010010001101100010011000001001111100000011011000000010111001111001001000010001010100110000000110110010001100011111000100101010001011010000100010000010000000000001101100000000000101000000000100),
      .INIT_6(256'b1100000001110011110110110101000111001000110100110101001101011001111010100101000111011011111110011100100001110111100001011110011011100010111110010100110101000000110000011000100110011111011110011110100110100011010010001000101011001000011100111101100111011001),
      .INIT_7(256'b1100100110000010100101011111011111100010111110010100100001010101010010001101001111001001011101110100100110000001100011000011110111000001101000001111001111101011010010010000000001011000110010101100000100100010110101011101110111001001100000100101110111001101),
      .INIT_8(256'b0110000011110100101100010010111111000000011100110101100101111011110010000111001110110000001110001100000001110011000010000110110111001001001000101000010010111001111000010010001001001100000000001100000110001000010010101101101101001001000000000100000100101010),
      .INIT_9(256'b0110100001010100010101101001010011100000010100111111100101111001111000000101001111111001011110011110000001010010110110010111110111001010110111001101001000000001111000000101001011111101011100010110101011110000110111010001100111000000110110110101010010011001),
      .INIT_A(256'b1110000110000010011111000101010101001001100010111001000101100011110010101110011011011101011001110100100011011001100101010011001111001010111001001101110001100010110010001111010110111010000100011100101110100011110010000110011111001011101000111110000001111001),
      .INIT_B(256'b0100000000111011000010001000011001100100110000010010110010000100110010101011000110000100001000101100000010011001100010100010001001101100111000111100000110100011010011100111111001001000000000000010010010000000001100010001101010011010000000010010010000000000),
      .INIT_C(256'b0100100011001100100000000110001000001100100011001101100100101001100011101010010011001001001000111111011111110101101100100100000101000100110001000000110010000110011011011000000110001010101000111100010000100010100001001000110111001010001110010010110010100011),
      .INIT_D(256'b1010010000101100110001000011001100000000000101101111100110000010111000000110110011011000011000111000111010100111110001000011100100001100100011111101010000110110000010001000111011011001001010001000111010100110110111000011011010001110101001001100000100101001),
      .INIT_E(256'b1010010000111000110000100001001111001010111001001001100000110011100111001101100110000110000000000100110000110011111110010110001011100000011010101101100101110110010111010010000010100100011000101010000000101111111101010010100000000100010111011101101001000001),
      .INIT_F(256'b1110000010010011011110001001010011001000100110010000010010101100010011001001001100100100100010000110000110001001011100001100100000100100100010000110000110000001011010010100000010100100001110011100001000010011100011101010001110011100001100111110000111000000)
    ) ram5 (
      .RDATA(memory_data_out_5),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1001010010011011110000110110000001001101010100000110101010011011100011000100110000111100000100011010101000011111111101110000000010101001011000100101111000000000100000000110101100001000100001101100111110101010100010010111011110000100111000011011110000100000),
      .INIT_1(256'b1011111000100111000001000010000011001111011000110100000000010001100001100111001101000100000100011110111101100010010000000001101110001110011100100100111010010001111000000100011110101101011011001011000001010010111011010111100111100000000100111010110001101101),
      .INIT_2(256'b0010001100101100010101010000100010101010010001000101010100000001010101110010001001000000011001001110001001010001000001011001110100001110000000000100010001000110000001001100011010010001000000010110000011010010000100010010010000100110000000000100000001010010),
      .INIT_3(256'b1010100001111001010100000100100111100010010100000001110010001101101011000010100001001000110011011100111000000110000100000101000010001100010100010100000010110001110001110100000101000100000110010010011001111000010000000001100101100111011010000100010000011001),
      .INIT_4(256'b1000010010100010100010001100111001011100010001001110101110001010101100100000000111010000111000010111011001011100010011010000000000011001110001011111101001000001110010101111100010011100001001110010110000000000000101000000000001010101100101100101100110001010),
      .INIT_5(256'b1011010000100010100010010110001000001000110110011101000001100011101001000111000111011100001101100000000010000110110110110000000010000100110110000101111010111100000011000101000011000101101000111000000010001000010011000000000001000010110110111111101000010001),
      .INIT_6(256'b1000010110001010011100100100100100100000101001000000100110001010100000010110001010000101110011001101101001101001110111011011011101011101100010001000010000100010110100001100100110001110011100101100110110100011011010000101000000011001100011101000010000100010),
      .INIT_7(256'b1100010111110010100010001001111001001101010100010100110010110110110001010111001001001100000100111100110101110011010010001011000011000101011100100100100000010000110110000010011011000001100010101100000001111010001101001010010110001110101010101001010000100010),
      .INIT_8(256'b0100110101010000001010000001010011001111111110011001010000110011010000000100011011001101110100101110000000110011110001010111001000011100100110111000100101100010111001010111000110000100001101100100110111011000100010000011011011101101110110111010111000010100),
      .INIT_9(256'b0100100000010001110001011101101100110110000110010110000111100000010011011101001011000000001100111100111111110010100111000011001100001000110101011000010001100011110010101111000010011001001001101000111010101000111011110101000111000000101100011000110011000110),
      .INIT_A(256'b0100110111010001100000000011001111000101111100000110011000011001010010000101010100101101010001001010110010001000111000100101000111000101111101001001101001011000010110010001000011000111000000100100101011010000000111000000010110000110000000100100111111011011),
      .INIT_B(256'b1100111010110011100010010010011011010101101000101100101011111001010011000100010110000100101010100000111011011001010010000001000100101100000000010100110010010001000001000111001001001000100100111000010000100010110001001011000100110010010010000101110100000000),
      .INIT_C(256'b0100010111100110101100100101000011110101010001011111100100100000111000000101001010010001001011000000010000000000100000100110001011100101100010001110010101010011110111000011100110001110111000011100110000110011110001011111001011110000001100110000110001000000),
      .INIT_D(256'b1000111010100010110000000111001001111100000100001010010000000010101111000010100001000101010100011001101000110011101011100110101101000110000100011000000000010000111110010000000011100101010100101001100000111001100001001100101001100110000110010110000011110000),
      .INIT_E(256'b0000110010100110110110001100001110010110000000000110111111111111010110000001010001000000110001000000011101000101000100000101001010001010001001111010010100000010110011010111110111010100101101101111111101101000001000011010000011001010111100011000010100111101),
      .INIT_F(256'b1000111010000010100001000010001001001100110010011100100011000111100110111000110010010000011100101101111110010000110100010010001001000010111110101001100110000110100001001010101001001010110110000101110000010000100001001010000011111101011001010101110100000000)
    ) ram6 (
      .RDATA(memory_data_out_6),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1010111000010101110101001100100101100001010010001110010011100110101000110000101011111110010000010100000011001100111001011100001011110110100111001010111101000000010001110101101111100100100100101110110111110010111011100001010001101111111011111110000010010011),
      .INIT_1(256'b0100000011100110110111011001001011001011101010101100010001100000000010001010010110011100011010010100001101101000111001100100010001011110010000001011110001000001010000001100110011100111010000011101000010011100011101010001001011100101101000100100010011000010),
      .INIT_2(256'b1111110111000100111010011000000000000000010001001001011001100011110001011110110111111010000101100111010110110100100000011010000011101000011000000101110101000001010001010010101010011100100100100101010011000001010011110100010011110100000101101010110101100000),
      .INIT_3(256'b0100110101010001100010101011000111000101011100111100010110110011111100100000111101001000000101001101010111101101111001000000011001001101010100011100101010011001101001100000000001000100111000111110010111010010111000000001000110000101001010001010000011001001),
      .INIT_4(256'b1101010001100010110100001010110111001100100111100100100001010000010101001001000010000100101000001100110111010011000010000001000111000111010100110100001000110000000011010000000001101100000000001000101011100011110101010010001010000100101000101111001001001011),
      .INIT_5(256'b0100000010011011101001100000000101001100100100010000010001010000110010000001100110001110001010101100010000110011100110101110001010001100011100101100111000111001100100000110001010001110111100011100110000110011100111101000001011010100011010001101101110000000),
      .INIT_6(256'b0000110101000000000011001101001011000100001100010100100011010100110000010110000110101110100010001010001000000101110101011010000001100010010111000100100101000001101001001000100010100100100110011110010010011100100001001011001011001100100110110000110001010001),
      .INIT_7(256'b1110011000010001000011001110000011100110000101101010010111010001111111011000000011101000110100011110110011000101101011001000000000010010000001101110111100000000010011011011010111110110000100110000010011110011110011001001001111000111000101100101011000110001),
      .INIT_8(256'b1001000100100110100011101000001010001100011100101100111110100000110000000110011010001111110101001000110000100010010010001101001011010100001100101000111000101010100011000010001001001100110000011100000001110011110110110111110010001100001000101010111011001001),
      .INIT_9(256'b1111110011000010000010001010101111011001001000101100111110010100110101000011011001001101101111000110100000110011010010001101011000010110010100010011100011111000111010100101010011010000100010010000010000000000110111010000010101010011100000001100101011110010),
      .INIT_A(256'b1010010101100010000011001111101111001100001101100000010001111000111001100001000101001000011100001110110001100001000011001010100010001001011010001101111110000000110000100000001001011000101010001101101000000011110011101001001011000101001101110100000000010100),
      .INIT_B(256'b1000111011010011111010000011100110111100011000101010011001010000110010101001000110111100011010000100100110101011111010000011110000010000010110001010011001010000010010001011100111010000011011001010100010000001011001011000100010101010000001000101110001100011),
      .INIT_C(256'b1100100000110011000111011111111110000100011000111100101011000110100100000010011101001100011100110110100001100110100001111100010100001100101010001000000001110011110011101100000111010101011001110000110100100000011011010111011111101100000100111011011000000000),
      .INIT_D(256'b0100110001110000110010110000001111000001110111110011001001011000001000001110010001001100110010011111010101101001010100010010001011000111010101011111000000111110111010010010001101001100101011101000110000100010101000000011110111111101001000100100110111111101),
      .INIT_E(256'b0100110111111110101001000010100000000100010110011110001000010000010110001010100011001000001110010000110001110000111000000011100100001101001000101110010001101001000000000100110111100111000000000100110101110101110010000011100001001000111011001001001000010010),
      .INIT_F(256'b1101010100100011110111111000000010011101011101111010110001000011111100100000000011001110101101101010100000100000010011001010101011001000011011001010110101101010101001100000000011001010101000001110100000110001010010001010100010010000001110011110000011011001)
    ) ram7 (
      .RDATA(memory_data_out_7),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b1101100001100010010011011111100011000001001000110000110011100000110011000011001100000001100101111111011100000000000001000100001110001010001100110000010011100010110011100001000110000100000100011110000010010011010001010100000111001110001100110000110010111000),
      .INIT_1(256'b0000110011101010110011010111000001001001101000111100110100110110010011001011100010000000011000100100100011110000100100010010010000001100101010001100110100110100010010001011000011011000011000100110110101010000010010011010101110000100011000110100110010110011),
      .INIT_2(256'b0101110101010101110011101110001110000000001001100101110110000010110010000010001010001110111000011000000000100111010011011001000111001000011001110110100100000100000001000000000011001000010001010000100011101110100100000111001001011101101001101101000100100000),
      .INIT_3(256'b0001110001000000100010101010010111000001001100111010000000101101100111110001001100111000010000000001110001101010100000000010011011100001001110111000100000100110000111010011100110010000011000101110010101111001110010000011001111000101110110101110001010011001),
      .INIT_4(256'b1111000100101000101000000010001100001001000110011000100000100010111001010011101110101001001010010100010000001000111000110000000011100000001010011010110000101000100010101010011110000001001000101110010101101101110010100001001110000010000000110011000100111001),
      .INIT_5(256'b0011000010110001100100101100000010001010101000011101010100110011110001110101001101101100000110010001100001000000100000001000101001110111000110010110010111110000111011000011000110001111010000001110000001101111101110010010011000011000010110101000100000100111),
      .INIT_6(256'b1000101101101010100101000110001010011110111000101100100100100010100101011010101000011010110110000000110101000000110011110111100011000000001100111001111011100000110011010111001111000000101110110001111011001000000010000100010010000101101000101110010101010001),
      .INIT_7(256'b1100011000010110100000000101000100001001000000000100010101000101110011101011000101111001111000010101001110000000110010100110100011001101011100111000111000111110110011010111100010000100101111100000101010001101000011010001010010001010101001001000110100110100),
      .INIT_8(256'b1100100100000000100111111111010110000100001000000001010000001000100010000000000101101001000100010000000000000001111111010001000101001001111000101000000000101000110000011011001110100000001000100111010110110001110000011110001000001111011010100101100000000001),
      .INIT_9(256'b0001110000000000001010000000010111000011000100010010000010000111001101011011000100000000000010111110011100010001000000001000010011100001100100111000101010100100100111110001001100000000000000001100110100010001110010101110011111000001001001000000110010000010),
      .INIT_A(256'b0000111110111100000010000010010010000001100111000100111111011011011000001011000100000000000001011100110110010011010001010101100001001010000100011000000010001100011001010001101100001001101000001110111010101010110010001100011111000001100011000000111010001010),
      .INIT_B(256'b1000100000000101111001110011000100100000001001100110000110110001100000001000101000011101101100010000001000000110010001110001000100100011011010000000100011011001111000010010001001100111110100111010110000010110010001110101000000001100001111101000001000000111),
      .INIT_C(256'b1010100000000001110011111011000000001010000000001110010110111011011001100110010011000000110100011111000110101111001001000010101010010110001000000101011010110110010100110000101011101000010000001000101010100101010010110001000110001010101000111001010100010001),
      .INIT_D(256'b1000000000001011111001110001100101100010010001011100001100010000000001100010100000010111011100011110110000000100110010101111000101011010000100011011000001011000001000100010001001100011000110101101000000000001010001100011110001010010000000110101001000010100),
      .INIT_E(256'b1000110010100000100101000000101000101000101010110110001110010001000111000100001010001000000010001100000110111011000101101110001011101100010001101100101011011011110100011000010100101110000000101011100001100010101000100010000001100101101110010011000011000010),
      .INIT_F(256'b1110010000101100001000001000011011010011000000100010010011010000010011000000010010011110101000000000111001000101010000101011001101001101010110111110110000010001100001100100111001001000001100011100111111011000110001000001101101100011001000110000110101001101)
    ) ram8 (
      .RDATA(memory_data_out_8),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0100100101000100000010000101000100001101010000000000100101010001000010010101000001011000010101000001100000010001000110000100000000010001000100000100000000010000010001010101000000001101101010100000010100110000000001011000001101001101111110101000011100100010),
      .INIT_1(256'b0100101000101001000110010100000101111100101010010010110010111111011010110000100100101110001000000010110101011111001011000011001001111110001111010000100100000000010011000000000001011001000100000001100100010001000110010000000000011000010101000001100001000001),
      .INIT_2(256'b0001000100000100000100010001000100010001000100000001000000010001000100010000010001000000010000010000000101010001111111101010101000010000111100110110110001011010011010001000011000101011000010110010100100000111011011010101100000001101000000000100111001110010),
      .INIT_3(256'b0101010001010000010100010001000000010001000001010001000001000001000100000101000001000001010000000000010001010001010101000000000001010000000100000001000001010100000100000001000101000000000100010000000101010001000000010001000101010100000000000101000001010100),
      .INIT_4(256'b0001000100000000010101000000000101000101010100000000010100000000000000010101000100000100000001010100000100000101000001000001000000000001010101010100000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000010000010000),
      .INIT_5(256'b0000010001000101010100010000010000010000000000010001000000010001000100000101000000010000000001010100000000010100000000000100010000000101010000000101000001010100000100010001000100010001000001000100000000010001000100010100000101000100010100000100000000000000),
      .INIT_6(256'b0001010000010000000000010001010101010001000001010000010100000000010001000101000101000000000100010000000100010000000001010100000001000101010100010100000000000000010001000000000000000001010100010101000001010001000100000001000100010001000001000100000000010000),
      .INIT_7(256'b0001000100010000000000010100000101010001000001010000010100000000010001000101000101000000000100010001000101000100000000010100000001010001000001010000010100000000010001000100010101000000000100010101000100000101000001010000000001000100010001010100000000000001),
      .INIT_8(256'b0000010001010101000100010001000000000001010001010101010000000100000001010000000001000100010101010100000000010001000100010100010000000001010001000101010000000100000001010000000001000100010001000100000000010001010101000000010000000101000000000000010001010101),
      .INIT_9(256'b0000000101000000010000000001000100000001010001000000000001000100000000010100010000000100010000010000000001000001000000000100010000000001000001000100000000000000010000000000000000000000010001000101000000010000000100000101010000010001000001000100000101000000),
      .INIT_A(256'b0000000000000101000000000001000100000000000001010000000000000100000000000001000000000000010001010001010100000100000101000000000100000101000000000000010100000001000000000100010100000000000000010000000100000100010000000000000000000000010000010000000100000101),
      .INIT_B(256'b0101000100000100000100010000010100010001000100010100000001010101000001000101010100000001000101010000000101010000000000000000000000000000000000000000000001000100000000000001010000000000010000010000000001000101000000010100000100000001010001000000000101000101),
      .INIT_C(256'b0101000000000001000001000101010100000001000001000100010000000100000001000101010100000100010101000100010001000001010000000000000000000100010001000000010100000001000001000100010000000101000000010100010101010000000001010000000001000100010000000100000000000000),
      .INIT_D(256'b0100010001000000010000000000000000000100010101010000000001000101010001010101000000000101010000000100010001010000010000000000010100000100010101010100010001000001010000000000000001000101010100000000010100000000010001000100000001000000000000000000010001010101),
      .INIT_E(256'b0100010101010100010000000001000000000100010101010100000100000101000000000100000101000101010100010100000000010000010001010101000001000000010101000000010001010101000000000000010000000000010000010100010101010001010000000001000000000100010101010001000100000100),
      .INIT_F(256'b0000000001000001010001010101000001000000000100000000010001010101000000000001010000000000010000010100010101010001010000000001000001000101010101000100000000000000000001000101010101000001000000010000000001000001000001000101010100000000000100010000000001000001)
    ) ram9 (
      .RDATA(memory_data_out_9),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram10 (
      .RDATA(memory_data_out_10),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram11 (
      .RDATA(memory_data_out_11),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram12 (
      .RDATA(memory_data_out_12),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram13 (
      .RDATA(memory_data_out_13),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram14 (
      .RDATA(memory_data_out_14),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram15 (
      .RDATA(memory_data_out_15),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram16 (
      .RDATA(memory_data_out_16),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram17 (
      .RDATA(memory_data_out_17),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram18 (
      .RDATA(memory_data_out_18),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram19 (
      .RDATA(memory_data_out_19),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram20 (
      .RDATA(memory_data_out_20),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram21 (
      .RDATA(memory_data_out_21),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram22 (
      .RDATA(memory_data_out_22),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    SB_RAM40_4K #(
      .READ_MODE(1),     // 512x8
      .WRITE_MODE(1),    // 512x8
      .INIT_0(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_8(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_9(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_C(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_D(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram23 (
      .RDATA(memory_data_out_23),
      .RADDR(rom_address),
      .WADDR(0),
      .WDATA(0),
      .RCLKE(1'b1),
      .RCLK(clk_40mhz),
      .RE(1'b1),
      .WCLKE(1'b0),
      .WCLK(clk_40mhz),
      .WE(1'b0)
    );

    ////
    // END - BRAM insertions.
    ////

endmodule
